module JK_flipflop (q, q_bar, j,k, clk, reset);
input j,k,clk, reset;
output reg q;
output q_bar;
// always@(posedge clk or negedge reset) // for asynchronous reset
always@(posedge clk) begin // for synchronous reset if reset)
  if (!reset)
    q<=0;
else
begin
case({j,k})
2'600: q < q; // No change
2'b01: q <= 1'b0; // reset
2'b10: q <= 1'bl; // set
2'b11: q <= ~q; // Toggle 
endcase
end
end
assign q_bar = ~q;
endmodule
